// DSCH 3.5
// 5/10/2023 7:28:35 PM
// example

module example( );
endmodule

// Simulation parameters in Verilog Format

// Simulation parameters
