// DSCH 3.5
// 5/11/2023 4:49:17 PM
// C:\Users\stanl\Documents\Univeristy\vlsi\dsch3.5\MUX_2_1.sch

module MUX_2_1( );
 wire w2,w3,w4,w5;
 mux #(1) mux_1(w5,w2,w3,w4);
endmodule

// Simulation parameters in Verilog Format

// Simulation parameters
